import uvm_pkg::*;
module test();
    initial begin
        run_test();
    end
endmodule